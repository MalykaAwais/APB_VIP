package apb_pkg;

 import uvm_pkg::*;
 `include "uvm_macros.svh"
  import param_pkg::*;
  typedef uvm_config_db#(virtual apb_if) apb_vif_config;

  `include "apb_master_packet.sv"

  `include "apb_master_monitor.sv"
  `include "apb_master_sequencer.sv"
  `include "apb_master_driver.sv"
  `include "apb_master_agent.sv"
  `include "apb_master_sequence.sv"

  `include "apb_master_env.sv"

endpackage : apb_pkg
